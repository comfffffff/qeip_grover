
`define USE_SRAM
`define SRAM_HEX_SIZE 7446
`define CRM_HEX_SIZE 0
`define DRAM_HEX_SIZE 0
`define HEX_SIZE 7446